// SOPC.sv
// Minimal SOPC