// MEM_WB.sv
// MEMory Phase to Write Back Phase