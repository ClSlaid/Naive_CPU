// EX_MEM.sv
// From EXecute Phase to MEMory Phase.