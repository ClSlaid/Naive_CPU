//ID_EX.sv
// EXecute phase