// naive cpu
// author: ClSlaid <cailue@bupt.edu.cn>

module Naive_CPU();
	if_pc pc0();
endmodule
