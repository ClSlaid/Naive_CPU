// ROM.sv
// Read Only Memory
