// mem.sv
// operation in MEMory Phase