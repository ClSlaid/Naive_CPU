// ex_alu.sv
// 