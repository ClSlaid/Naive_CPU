//de_unpacker.sv
//author: ClSlaid <cailue@bupt.edu.cn>
